`define RF_PATH   CPU.EXstage1.RegFile1.rf
`define DMEM_PATH CPU.EXstage1.DMEM1.dmem
`define IMEM_PATH CPU.IFstage1.IMEM1.imem

